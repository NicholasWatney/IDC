

module test;

    reg clock;
    reg [15:0] A;
    reg [15:0] B;

endmodule

module adder(
    input clock,
    input [15:0] A,
    input [15:0] B
    );

    wire clock;
    wire [15:0] A;
    wire [15:0] B;

endmodule
